library verilog;
use verilog.vl_types.all;
entity Arithmetic_LU_vlg_vec_tst is
end Arithmetic_LU_vlg_vec_tst;
